LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY random_rom IS
PORT (
      clk          : IN  STD_LOGIC;
      address         : IN  STD_LOGIC_VECTOR(9 DOWNTO 0);
      random_value       : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
      );
END  random_rom;

ARCHITECTURE Behavioral OF random_rom IS

  TYPE rom_type IS ARRAY (0 TO 999) OF std_logic_vector (7 DOWNTO 0);
  SIGNAL memory : rom_type :=(
  "01010000","01011000","10100100","01000001","01110100","00110001","01011010","01100011","10100000","10011010","00110101","01100100","00111000","10000000","10000000","01101101","01111100","10000011","10001000","01100111","10100011","00110101","10010100","10010101","01100011","00111001","01100010","10010011","10011101","01010000","01111011","10011110","10000001","10011100","01001010","10001011","10001000","10000101","01010110","01110000","10011110","01100110","00110111","01011100","00111011","01100100","00101010","01101111","01110011","10010100","01100011","10001000","01101111","00110011","01001101","00111010","01000101","00110001","01011001","00111000","01110100","10000000","01000000","00111011","10010101","01111111","00101001","00111110","10011101","01001111","10001001","01010010","01010011","00101110","01100011","01011100","01111000","01000001","01101010","01000011","10010111","10001110","01100101","10011100","00101111","00110011","00110110","01001110","01100000","10000111","01110010","10010111","01101010","00101001","01101011","00111000","01011110","01001010","01100011","00101100","01100111","00111000","01010011","00110110","00111010","01110101","01101110","01110101","01010101","01100000","00111101","10011001","10011111","01110111","10010011","01001000","01010110","00110010","10100100","10000100","01110010","01101011","00100110","01001101","10011010","01101000","01000101","01001110","10100001","01001100","01110001","01000110","10001000","01011010","00110101","01101110","01001010","01101101","10010111","00111110","00111011","00101110","01001001","01100101","01010110","10001111","10001111","01111000","10011011","01001001","00111001","10001001","10011000","01010001","10010011","01100011","01100111","01001000","01000000","01110001","01101101","10001100","00111011","01000101","10100000","00101010","00110111","01101010","00101110","01010001","01001111","00110000","00100110","10011000","10000000","01011101","10001001","00110110","01100011","10000011","01111110","01111001","01100001","01101011","10010000","01000100","01001010","10010111","00110110","01100110","01010001","00111001","00110010","01000101","01001111","01101001","10001011","10011000","01100110","00101010","01000100","01000010","00111010","01010100","01101100","01100011","10000111","10011100","10010000","01010110","00111110","01010001","10011001","10100100","00111001","00110001","01101010","01010100","01100000","10001100","00110111","00100100","10011000","01000001","10100010","01001101","10001100","01001000","10011100","01110100","10001100","01100100","10000010","10001010","00110111","01000100","01111101","01110110","00101011","10011110","10011100","00101001","01111100","10000111","01010111","01010110","00101111","01111000","01101111","01001101","10011010","10100010","01110100","00101111","01010100","01111111","01111101","00110100","01110011","01010001","00110100","01110010","01101101","10001110","01011011","00100110","10001001","01001001","01111001","10010001","01011000","10000100","00100011","00111101","01000100","10100001","10100010","01111110","00111101","01010000","00101011","00101000","10011100","10011011","01110001","10011110","00110011","10000001","00110011","01011011","10001111","00111001","01000100","01100001","10000000","01000100","01000110","01110111","01000110","10000110","10011001","10011000","00111011","10000111","01001110","10001100","10010000","10010010","01010100","00110111","00110011","00100111","10000111","00101000","01011001","01010010","00100100","00111100","00111000","01001010","01000101","10001111","01110111","01011101","00101111","10010110","00100100","01111011","01000010","10010010","01101001","10001010","01101001","10011111","01010010","01111010","10011000","01100000","00110111","10100100","01101000","01111011","01100101","00111001","01101100","00110111","01010010","10000000","01000000","01011101","01110111","10100000","10000101","00110000","10010010","01000111","10010011","01111001","00111010","00101001","00101011","01100101","01100011","10100010","00100101","10100001","10011001","10011111","00110111","01111000","00101100","10000011","01101010","01010111","01110010","00101001","01111110","10011000","01100001","01001000","10000011","01111011","01001101","01001100","01001111","01000101","10011000","01000100","10010100","10000100","10001011","01110101","10100001","01011110","01000001","01110101","01011111","01111101","01001000","01110000","01111001","01001110","00110100","01000110","01110101","01011010","01001111","10000101","00111110","00100100","10100010","10000110","00110101","00100100","01100101","00101001","10010111","01101001","01100100","00110011","01100000","01000000","10000010","01110000","00110011","01011011","10000001","01100101","10000111","10001101","00101100","10001101","00111011","00111011","00111000","01001010","10010011","01001111","01111100","00110010","00110011","10010100","01010110","00100100","01100111","00100110","01011111","10010000","01010100","01001010","10100100","01001101","01011010","01010000","01101000","01011101","01111101","01100000","01101011","01011001","01000111","00111101","01101111","01101111","10010000","00101100","00100111","01001111","01010110","01100111","00101000","10000110","01000000","01010100","10100000","01100011","10001001","01011101","10001010","01001010","01110111","10011100","01010010","01111011","00110100","01001010","01100101","01111110","00111110","01111111","01100000","00110011","01011000","01111001","10011000","01111010","01100100","01001001","10000101","10011110","10100011","01110000","01001110","10010001","10000100","01101001","01011100","01011101","01001101","01001111","10000001","01101110","01101010","10011110","01101001","00110010","10011001","00100110","01111001","10010010","01100100","00111100","01110101","01010110","00100111","10000100","01100111","10000111","01111010","01010110","00110000","00101100","01011001","01011101","00110010","10011100","01011011","01010100","10100000","00101011","01110011","00101000","10010000","10001011","01111001","00111110","00111110","00111000","01011000","01101100","01110101","10000101","01010010","10001101","01001101","10000100","00110111","01100001","00100101","10010100","01001010","01010111","10011110","01110010","01110111","00110010","00111101","10001110","10011101","01010010","10001110","01001001","01011000","00111011","10011100","01011110","01010100","10011101","00101001","10010001","10011001","01101010","01111001","10001101","10010000","01011010","01111010","01011110","01001000","01001101","01001110","01010010","10000100","10100100","10000001","00100011","01011100","01011110","00110100","01111010","01001000","01100000","01100101","01000001","01010010","10010010","10001111","10000000","10000101","01011100","01100011","00101010","00110011","01010000","01010000","01001000","10010110","01000000","01001011","01101010","01100001","10000110","01000000","01011100","01010010","01010101","01100110","00110011","10010100","10011110","01111001","01100110","10100011","00101111","00111110","00111000","00111101","01110100","01101000","10010010","00110010","10100100","10010010","01000101","01001110","01111111","10011101","01110011","10001010","10011101","00101011","00110101","01000110","10001001","10011111","01000110","01110101","01100101","01111010","00110001","00100100","01010111","10000000","01001110","00110101","01001000","00111110","01111100","10011000","01110101","10100001","01111011","01011010","01101011","01111101","10001110","00101101","00110001","01001110","00110110","01000101","00100110","01100010","10000110","00100100","00111000","01110110","10011111","01000000","01010011","01110110","10100000","01110001","01100001","10010100","01001100","00111000","01111111","00100101","01101010","00101110","01111101","10001001","01001110","01100001","00110100","10010100","01000101","01101000","01100011","00101110","01100011","01001011","10000101","10000011","10100000","00101111","01100000","01110110","00111011","10010111","01010001","00100100","00110001","00110011","01010111","00101111","00111010","01100011","10100100","01110100","01011111","10000010","00101011","01110010","01011101","01100100","00111100","01100010","01011110","00111010","10011111","01011000","00111111","10010010","01111011","01110100","01101110","00100011","00110001","10000101","10000000","01111111","10010111","01110011","00110111","00111100","10000001","10010101","10000100","01111111","01010000","10100001","00110110","01100001","00101100","10001000","10001110","10011010","01001011","00110100","00111110","10011100","10001011","00110001","10011111","10010001","00100011","01101100","00110101","01001111","00111111","10001100","10010101","01110111","01100110","00111010","01101100","01010101","10010111","10000100","00110100","01110000","10010011","10011001","01101100","00101000","01010100","00100110","01011110","00110010","01101000","10001001","00101010","01011110","10011111","01111000","01011010","00111100","00101101","00100101","01001000","01110111","01000010","10011001","01101101","01101100","10000000","10000110","10001011","10001000","10010111","01111100","00101010","00110100","00110001","00110010","10010000","01011100","10010000","00101000","01010011","01110000","01110100","01001101","01010011","01000110","01001110","01001010","00110001","10000011","01100111","01000110","10011001","10011111","01001001","01101000","10010010","01010101","01010101","01101001","01101101","01110000","01101100","01101101","10010011","00110101","01110101","10011010","00111001","10000001","10001111","01011001","01100011","01000101","10011000","10010000","01000010","00111101","01010000","00101110","01010110","10100001","10100100","10001110","10011010","00111101","01010101","01100000","10000011","01110000","01101100","10010100","01110000","01101101","01001010","10100011","10000011","10001000","01110011","01100010","10001011","01011110","00111001","01000010","01110111","00101010","00111011","10000100","01011010","10010010","10001000","01010101","00101111","10000110","10011101","00110101","01011100","10010111","10010111","01111001","00101100","01101110","00100101","01100101","10010010","00110101","01000010","10011000","10000001","10010001","00110110","01000111","01111110","01111111","01000110","01001110","01010110","01010100","00100110","10001101","01010100","10011100","00101110","01000010","10010110","10100011","10011000","01010010","01100000","00101110","01111011","00110001","00110111","00101110","10011100","00100011","10011011","01100010","10000001","00100100","01010010","01000010","10011110","10000001","01001100","01011110","10000111","01011000","01101101","10010100","01010011","00101011","00101111","10010000","10100011","10010010","01000100","10000011","01100011","10100010","10010010","10100011","00110001","01101100","00101101","10011000","01110011","10001010","10011101","10100001","10011011","01000110","10010110","00110111","10010101","10100000","10010001","01110001","10001000","00100110","01110100","00110111","01000000","01011111","01111111","01101000","00100100","01101000","01011010");
      ATTRIBUTE RAM_STYLE : string;
  ATTRIBUTE RAM_STYLE of memory: signal is "BLOCK";

BEGIN

  PROCESS (clk)
  BEGIN
    IF (rising_edge(clk)) THEN
      random_value <= memory(to_integer(UNSIGNED(address))) ;
    END IF;
  END PROCESS;
  
END Behavioral;