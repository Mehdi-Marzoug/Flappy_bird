LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY game_over IS
PORT (
      clk          : IN  STD_LOGIC;
      address         : IN  STD_LOGIC_VECTOR(12 DOWNTO 0);
      pixel_game_over       : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
      );
END game_over;

ARCHITECTURE Behavioral OF game_over IS

  TYPE rom_type IS ARRAY (0 TO 4999) OF std_logic_vector (2 DOWNTO 0);
  SIGNAL memory : rom_type :=(
  "111","111","111","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","100","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","100","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","110","110","110","110","110","110","110","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","000","111","111","111","110","110","110","110","111","111","111","100","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","110","110","110","110","110","110","110","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","100","000","000","000","000","000","111","111","111","111","111","111","111","111","111","000","111","111","110","110","110","110","110","110","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","100","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","110","110","110","110","110","110","110","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","100","111","111","111","110","110","110","110","110","110","111","111","111","100","111","111","111","111","111","111","111","111","111","100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","110","110","110","110","110","110","110","110","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","000","111","111","110","110","110","110","110","110","110","111","111","111","000","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","110","110","110","110","110","110","110","110","111","111","000","000","000","000","000","000","000","000","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","100","100","000","111","111","111","110","110","111","110","111","111","111","111","111","111","111","111","111","111","000","111","111","110","110","110","110","110","110","110","110","111","111","000","000","000","000","000","000","000","000","000","100","111","111","111","110","111","111","110","111","111","111","111","111","000","000","000","000","100","000","000","000","000","000","111","110","110","110","110","110","110","110","110","110","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","110","110","110","110","110","111","111","000","111","111","111","111","111","111","000","111","111","110","110","110","110","110","110","110","110","111","111","000","000","000","000","000","000","000","000","000","000","111","111","110","110","110","110","110","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","111","110","110","110","110","110","110","110","110","110","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","111","111","111","110","110","110","110","110","111","111","000","111","111","111","111","111","111","000","111","111","110","110","110","110","110","110","110","110","111","111","000","111","111","111","111","111","111","111","111","111","111","111","110","110","110","110","110","111","111","111","000","111","111","111","111","111","111","111","111","000","000","000","111","110","110","110","110","100","100","100","100","100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","110","110","110","110","110","110","110","111","000","111","111","111","111","111","111","000","111","111","110","110","110","110","110","110","110","110","111","111","111","111","111","111","111","111","111","111","111","111","111","110","110","110","110","110","110","110","111","111","000","111","111","111","111","111","111","111","111","111","000","000","111","110","110","110","110","110","100","100","100","100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","110","110","110","110","110","110","110","111","100","111","111","111","111","111","111","000","111","111","110","110","110","110","110","110","110","110","111","111","111","111","111","111","111","111","111","111","111","111","111","110","110","110","110","110","110","110","111","111","000","111","111","111","111","111","111","111","111","111","000","000","111","110","110","110","110","111","111","111","111","111","111","111","111","111","110","110","110","110","110","110","111","111","110","110","110","110","110","110","110","110","110","110","110","110","110","111","111","111","111","111","110","110","110","110","110","110","110","111","111","000","111","111","111","111","111","000","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","111","110","110","110","110","110","110","110","111","111","111","111","111","110","110","110","110","110","111","111","000","000","111","110","110","110","110","111","111","111","111","111","111","111","111","111","110","110","110","110","110","110","110","111","110","110","110","110","110","110","110","110","110","110","110","110","110","111","111","111","111","111","110","110","110","110","110","110","110","111","111","000","111","111","111","111","111","000","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","111","110","110","110","110","110","110","110","111","111","111","111","111","110","110","110","110","110","110","111","000","000","111","110","110","110","110","111","111","111","111","111","111","111","111","110","110","110","110","110","110","110","110","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","111","111","111","110","110","110","110","110","110","110","110","111","111","000","111","111","111","111","111","000","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","111","110","110","110","110","110","110","110","110","111","111","111","110","110","110","110","110","110","110","111","000","000","111","110","110","110","110","111","111","111","111","111","111","111","111","110","110","110","110","110","110","110","110","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","111","111","111","110","110","110","110","110","110","110","110","110","111","000","111","111","111","111","111","000","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","110","110","110","110","110","111","111","111","110","110","110","110","110","110","110","111","000","000","111","110","110","110","110","111","111","111","111","111","111","111","111","110","110","110","110","110","110","110","110","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","111","111","111","110","110","110","110","110","110","110","110","110","111","000","111","111","111","111","111","000","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","110","110","110","110","110","111","111","111","110","110","110","110","110","110","110","111","000","000","111","110","110","110","110","111","111","110","110","110","111","111","111","110","110","110","110","110","110","110","110","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","111","111","111","110","110","110","110","110","110","110","110","110","111","000","111","111","111","111","111","000","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","100","110","110","110","110","111","111","111","110","110","110","110","110","110","110","111","000","000","111","110","110","110","110","111","111","110","110","110","111","111","111","110","110","110","110","110","110","110","110","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","111","111","111","110","110","110","110","110","110","110","110","110","111","000","111","111","111","111","111","000","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","100","110","110","110","110","111","111","111","110","110","110","110","110","110","110","111","000","000","111","110","110","110","110","111","111","110","110","110","111","111","110","110","110","110","110","110","110","110","110","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","000","111","111","111","111","111","000","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","110","110","110","110","110","111","111","110","110","110","110","110","110","110","110","111","000","000","111","110","110","110","110","111","111","110","110","110","111","111","110","110","110","110","110","110","110","110","110","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","000","111","111","111","111","111","000","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","111","111","110","110","110","111","111","110","110","110","110","110","110","110","110","111","000","000","111","110","110","110","110","111","111","110","110","110","111","111","110","110","110","110","110","110","110","110","110","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","000","111","111","111","111","111","000","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","111","111","110","110","110","111","111","110","110","110","110","110","110","110","110","111","000","000","111","110","110","110","110","111","111","110","110","110","111","111","110","110","110","110","100","110","110","110","110","111","110","110","110","110","100","110","110","110","110","110","100","110","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","000","111","111","111","111","111","000","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","111","111","110","110","110","111","111","110","110","110","110","100","100","100","110","111","000","000","111","110","110","110","110","111","111","110","110","110","111","111","110","110","110","110","110","110","110","110","110","111","110","110","110","110","100","110","110","110","110","110","100","110","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","000","111","111","111","111","111","000","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","111","111","110","110","110","111","111","110","110","110","110","100","100","100","110","111","000","000","111","110","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","110","111","110","110","110","110","111","111","110","110","110","110","110","110","110","110","110","111","000","111","111","111","111","111","000","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","111","111","111","111","000","000","111","110","110","110","110","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","110","111","111","110","110","110","111","111","110","110","110","110","100","110","110","110","110","111","000","111","111","111","111","111","000","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","111","111","110","110","110","111","111","110","110","110","111","111","111","111","111","111","000","000","111","110","110","110","110","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","110","111","111","110","110","110","111","111","110","110","110","110","110","110","110","110","110","111","000","111","111","111","111","111","000","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","111","111","110","110","110","111","111","111","111","111","111","000","000","111","110","110","110","110","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","110","111","111","110","110","110","111","111","110","110","110","110","110","110","110","110","110","111","000","111","111","111","111","111","000","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","110","110","110","110","110","111","111","110","110","110","111","111","000","000","000","000","000","000","111","110","110","110","110","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","110","111","111","110","110","110","111","111","110","110","110","110","110","110","110","110","110","111","000","111","111","111","111","111","000","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","110","110","110","110","110","111","111","110","110","110","111","111","000","000","000","000","000","000","111","110","110","110","110","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","110","111","111","110","110","110","111","111","110","110","110","110","110","110","110","110","110","111","000","111","111","111","111","111","000","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","110","110","110","110","110","111","111","110","110","110","111","111","000","111","111","111","111","000","111","110","110","110","110","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","110","111","111","110","110","110","111","111","110","110","110","110","110","110","110","110","110","111","000","111","111","111","111","111","000","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","110","110","110","110","110","111","111","110","110","110","111","111","000","111","111","111","111","000","111","110","110","110","110","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","110","111","111","110","110","110","111","111","110","110","110","110","110","100","100","100","110","111","000","111","111","111","111","111","000","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","110","110","100","100","100","111","111","110","110","110","111","111","000","111","111","111","111","000","111","110","110","110","110","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","110","111","111","110","110","110","111","111","110","110","110","110","110","100","100","100","100","111","000","111","111","111","111","111","000","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","100","111","110","110","110","110","110","100","100","100","100","111","111","110","110","110","111","111","000","111","111","111","111","000","111","110","110","110","110","111","110","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","110","111","111","110","110","110","111","111","110","110","110","110","110","110","110","110","110","111","000","111","111","111","111","111","000","111","111","110","110","110","111","111","110","110","110","111","111","110","110","110","110","111","110","110","110","110","111","110","110","110","110","110","110","110","110","110","111","111","110","110","110","111","111","000","111","111","111","111","000","111","110","110","110","110","110","110","110","110","110","111","111","110","110","110","110","110","110","110","110","110","111","110","110","110","110","111","110","110","110","110","110","111","111","110","110","110","111","111","110","110","110","110","110","111","111","111","111","111","000","111","111","111","111","111","000","111","111","110","110","110","110","110","110","110","110","111","111","110","110","110","110","110","110","110","100","111","111","110","110","110","110","110","111","111","111","111","111","111","110","110","110","111","111","000","111","111","111","111","000","111","110","110","110","110","110","110","110","110","110","111","111","110","110","110","110","110","110","110","110","110","111","110","110","110","110","111","110","110","110","110","110","111","111","110","110","110","111","111","110","110","110","110","110","111","111","111","111","111","000","111","111","111","111","111","000","111","111","110","110","110","110","110","110","110","110","111","111","110","110","110","110","110","110","110","110","111","111","110","110","110","110","110","111","111","111","111","111","111","110","110","110","111","111","000","111","111","111","111","000","111","110","110","110","110","110","110","110","110","110","111","111","110","110","110","110","110","110","110","110","110","111","110","110","110","110","111","110","110","110","110","110","111","111","110","110","110","111","111","110","110","110","110","110","111","000","100","100","000","000","111","111","111","111","111","000","111","110","110","110","110","110","110","110","110","110","110","111","110","110","110","110","110","110","100","111","111","111","110","110","110","110","110","111","111","000","000","111","111","110","110","110","111","111","000","111","111","111","111","000","111","100","110","110","110","110","110","110","110","110","111","111","100","110","110","110","110","110","110","110","110","111","110","110","110","110","111","110","110","110","110","110","111","111","110","110","110","111","111","100","110","110","110","110","111","000","000","000","000","000","111","111","111","111","111","000","111","110","110","110","110","110","110","110","110","110","110","111","110","110","110","110","110","110","100","111","111","111","110","110","110","110","110","111","111","000","000","111","111","110","110","110","111","111","000","111","111","111","111","000","111","111","110","110","110","110","110","110","110","110","111","111","110","110","110","110","110","110","110","110","110","111","110","110","110","110","111","110","110","110","110","110","111","111","110","110","110","111","111","110","110","110","110","110","111","000","100","100","000","111","111","111","111","111","111","000","111","111","110","110","110","110","110","110","110","110","111","111","110","110","110","110","110","110","111","111","111","111","111","110","110","110","110","111","111","000","000","111","111","110","110","110","111","111","000","111","111","111","111","000","111","111","110","110","110","110","110","110","110","110","111","111","111","100","110","110","110","110","110","110","110","111","110","110","110","110","111","110","110","110","110","110","111","111","110","110","110","111","111","111","100","110","110","110","111","000","111","111","111","111","111","111","111","111","111","000","111","111","110","110","110","110","110","110","100","110","111","111","110","110","110","110","110","100","111","111","000","111","111","100","110","110","110","111","111","111","000","111","111","110","110","110","111","111","000","111","111","111","111","000","111","111","110","110","110","110","110","110","110","110","111","111","111","110","110","110","110","110","110","110","110","111","110","110","110","110","111","110","110","110","110","110","111","111","110","110","110","111","111","111","110","110","110","110","111","000","111","111","111","111","111","111","111","111","111","100","111","111","111","110","110","110","110","110","110","111","111","111","110","110","110","110","110","110","111","111","000","111","111","110","110","110","110","111","111","111","000","111","111","110","110","110","111","111","000","111","111","111","111","111","100","111","111","110","100","100","100","100","100","100","111","111","111","111","100","100","100","100","100","100","110","111","100","100","100","100","111","110","100","100","100","100","111","110","100","100","100","111","111","111","111","100","100","110","111","000","111","111","111","111","111","111","111","111","111","111","100","111","111","110","100","100","100","100","110","111","111","111","100","100","100","100","100","111","111","000","111","000","111","111","110","100","100","111","111","111","000","111","111","100","100","100","110","111","000","111","111","111","111","111","000","111","111","110","100","100","100","100","100","100","111","111","111","111","100","100","100","100","100","100","110","111","100","100","100","100","111","110","100","100","100","100","111","110","100","100","100","111","111","111","111","100","100","110","111","000","111","111","111","111","111","111","111","111","111","111","000","111","111","110","100","100","100","100","110","111","111","111","100","100","100","100","100","111","111","000","111","000","111","111","110","100","100","111","111","111","000","111","111","100","100","100","110","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","000","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","100","111","111","111","111","111","111","111","000","111","111","111","000","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","000","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","100","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","000","111","111","111","000","111","111","111","111","111","100","111","000","000","111","111","111","111","111","111","000","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","000","000","000","000","000","000","111","111","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","100","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","000","000","000","000","000","000","111","111","000","000","000","000","000","000","000","100","111","111","111","111");
    ATTRIBUTE RAM_STYLE : string;
  ATTRIBUTE RAM_STYLE of memory: signal is "BLOCK";

BEGIN

  PROCESS (clk)
  BEGIN
    IF (rising_edge(clk)) THEN
      pixel_game_over <= memory(to_integer(UNSIGNED(address))) ;
    END IF;
  END PROCESS;
  
END Behavioral;