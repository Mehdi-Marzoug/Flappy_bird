LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY pause IS
PORT (
      clk          : IN  STD_LOGIC;
      address         : IN  STD_LOGIC_VECTOR(12 DOWNTO 0);
      pixel_pause       : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
      );
END pause;

ARCHITECTURE Behavioral OF pause IS

  TYPE rom_type IS ARRAY (0 TO 2499) OF std_logic_vector (2 DOWNTO 0);
  SIGNAL memory : rom_type :=(
  "000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000");
    ATTRIBUTE RAM_STYLE : string;
  ATTRIBUTE RAM_STYLE of memory: signal is "BLOCK";

BEGIN

  PROCESS (clk)
  BEGIN
    IF (rising_edge(clk)) THEN
      pixel_pause <= memory(to_integer(UNSIGNED(address))) ;
    END IF;
  END PROCESS;
  
END Behavioral;